// traffic_light.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module traffic_light (
		input  wire       clk_clk,                          //                       clk.clk
		output wire [3:0] hex_0_external_connection_export, // hex_0_external_connection.export
		output wire [3:0] hex_1_external_connection_export, // hex_1_external_connection.export
		output wire [7:0] hex_2_external_connection_export, // hex_2_external_connection.export
		output wire [7:0] hex_3_external_connection_export, // hex_3_external_connection.export
		output wire [7:0] hex_4_external_connection_export, // hex_4_external_connection.export
		output wire [7:0] hex_5_external_connection_export, // hex_5_external_connection.export
		output wire       led_external_connection_export,   //   led_external_connection.export
		input  wire       reset_reset_n,                    //                     reset.reset_n
		output wire [2:0] tl_0_external_connection_export,  //  tl_0_external_connection.export
		output wire [2:0] tl_1_external_connection_export,  //  tl_1_external_connection.export
		output wire [2:0] tl_2_external_connection_export,  //  tl_2_external_connection.export
		output wire [2:0] tl_3_external_connection_export   //  tl_3_external_connection.export
	);

	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire  [18:0] cpu_data_master_address;                                   // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_data_master_read;                                      // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire         cpu_data_master_write;                                     // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [18:0] cpu_instruction_master_address;                            // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                               // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	wire         mm_interconnect_0_code_memory_s1_chipselect;               // mm_interconnect_0:CODE_MEMORY_s1_chipselect -> CODE_MEMORY:chipselect
	wire  [31:0] mm_interconnect_0_code_memory_s1_readdata;                 // CODE_MEMORY:readdata -> mm_interconnect_0:CODE_MEMORY_s1_readdata
	wire  [13:0] mm_interconnect_0_code_memory_s1_address;                  // mm_interconnect_0:CODE_MEMORY_s1_address -> CODE_MEMORY:address
	wire   [3:0] mm_interconnect_0_code_memory_s1_byteenable;               // mm_interconnect_0:CODE_MEMORY_s1_byteenable -> CODE_MEMORY:byteenable
	wire         mm_interconnect_0_code_memory_s1_write;                    // mm_interconnect_0:CODE_MEMORY_s1_write -> CODE_MEMORY:write
	wire  [31:0] mm_interconnect_0_code_memory_s1_writedata;                // mm_interconnect_0:CODE_MEMORY_s1_writedata -> CODE_MEMORY:writedata
	wire         mm_interconnect_0_code_memory_s1_clken;                    // mm_interconnect_0:CODE_MEMORY_s1_clken -> CODE_MEMORY:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;                   // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                     // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                      // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                        // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                    // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_tl_1_s1_chipselect;                      // mm_interconnect_0:TL_1_s1_chipselect -> TL_1:chipselect
	wire  [31:0] mm_interconnect_0_tl_1_s1_readdata;                        // TL_1:readdata -> mm_interconnect_0:TL_1_s1_readdata
	wire   [1:0] mm_interconnect_0_tl_1_s1_address;                         // mm_interconnect_0:TL_1_s1_address -> TL_1:address
	wire         mm_interconnect_0_tl_1_s1_write;                           // mm_interconnect_0:TL_1_s1_write -> TL_1:write_n
	wire  [31:0] mm_interconnect_0_tl_1_s1_writedata;                       // mm_interconnect_0:TL_1_s1_writedata -> TL_1:writedata
	wire         mm_interconnect_0_tl_0_s1_chipselect;                      // mm_interconnect_0:TL_0_s1_chipselect -> TL_0:chipselect
	wire  [31:0] mm_interconnect_0_tl_0_s1_readdata;                        // TL_0:readdata -> mm_interconnect_0:TL_0_s1_readdata
	wire   [1:0] mm_interconnect_0_tl_0_s1_address;                         // mm_interconnect_0:TL_0_s1_address -> TL_0:address
	wire         mm_interconnect_0_tl_0_s1_write;                           // mm_interconnect_0:TL_0_s1_write -> TL_0:write_n
	wire  [31:0] mm_interconnect_0_tl_0_s1_writedata;                       // mm_interconnect_0:TL_0_s1_writedata -> TL_0:writedata
	wire         mm_interconnect_0_tl_2_s1_chipselect;                      // mm_interconnect_0:TL_2_s1_chipselect -> TL_2:chipselect
	wire  [31:0] mm_interconnect_0_tl_2_s1_readdata;                        // TL_2:readdata -> mm_interconnect_0:TL_2_s1_readdata
	wire   [1:0] mm_interconnect_0_tl_2_s1_address;                         // mm_interconnect_0:TL_2_s1_address -> TL_2:address
	wire         mm_interconnect_0_tl_2_s1_write;                           // mm_interconnect_0:TL_2_s1_write -> TL_2:write_n
	wire  [31:0] mm_interconnect_0_tl_2_s1_writedata;                       // mm_interconnect_0:TL_2_s1_writedata -> TL_2:writedata
	wire         mm_interconnect_0_tl_3_s1_chipselect;                      // mm_interconnect_0:TL_3_s1_chipselect -> TL_3:chipselect
	wire  [31:0] mm_interconnect_0_tl_3_s1_readdata;                        // TL_3:readdata -> mm_interconnect_0:TL_3_s1_readdata
	wire   [1:0] mm_interconnect_0_tl_3_s1_address;                         // mm_interconnect_0:TL_3_s1_address -> TL_3:address
	wire         mm_interconnect_0_tl_3_s1_write;                           // mm_interconnect_0:TL_3_s1_write -> TL_3:write_n
	wire  [31:0] mm_interconnect_0_tl_3_s1_writedata;                       // mm_interconnect_0:TL_3_s1_writedata -> TL_3:writedata
	wire         mm_interconnect_0_hex_0_s1_chipselect;                     // mm_interconnect_0:HEX_0_s1_chipselect -> HEX_0:chipselect
	wire  [31:0] mm_interconnect_0_hex_0_s1_readdata;                       // HEX_0:readdata -> mm_interconnect_0:HEX_0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_0_s1_address;                        // mm_interconnect_0:HEX_0_s1_address -> HEX_0:address
	wire         mm_interconnect_0_hex_0_s1_write;                          // mm_interconnect_0:HEX_0_s1_write -> HEX_0:write_n
	wire  [31:0] mm_interconnect_0_hex_0_s1_writedata;                      // mm_interconnect_0:HEX_0_s1_writedata -> HEX_0:writedata
	wire         mm_interconnect_0_hex_1_s1_chipselect;                     // mm_interconnect_0:HEX_1_s1_chipselect -> HEX_1:chipselect
	wire  [31:0] mm_interconnect_0_hex_1_s1_readdata;                       // HEX_1:readdata -> mm_interconnect_0:HEX_1_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_1_s1_address;                        // mm_interconnect_0:HEX_1_s1_address -> HEX_1:address
	wire         mm_interconnect_0_hex_1_s1_write;                          // mm_interconnect_0:HEX_1_s1_write -> HEX_1:write_n
	wire  [31:0] mm_interconnect_0_hex_1_s1_writedata;                      // mm_interconnect_0:HEX_1_s1_writedata -> HEX_1:writedata
	wire         mm_interconnect_0_hex_2_s1_chipselect;                     // mm_interconnect_0:HEX_2_s1_chipselect -> HEX_2:chipselect
	wire  [31:0] mm_interconnect_0_hex_2_s1_readdata;                       // HEX_2:readdata -> mm_interconnect_0:HEX_2_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_2_s1_address;                        // mm_interconnect_0:HEX_2_s1_address -> HEX_2:address
	wire         mm_interconnect_0_hex_2_s1_write;                          // mm_interconnect_0:HEX_2_s1_write -> HEX_2:write_n
	wire  [31:0] mm_interconnect_0_hex_2_s1_writedata;                      // mm_interconnect_0:HEX_2_s1_writedata -> HEX_2:writedata
	wire         mm_interconnect_0_hex_3_s1_chipselect;                     // mm_interconnect_0:HEX_3_s1_chipselect -> HEX_3:chipselect
	wire  [31:0] mm_interconnect_0_hex_3_s1_readdata;                       // HEX_3:readdata -> mm_interconnect_0:HEX_3_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_3_s1_address;                        // mm_interconnect_0:HEX_3_s1_address -> HEX_3:address
	wire         mm_interconnect_0_hex_3_s1_write;                          // mm_interconnect_0:HEX_3_s1_write -> HEX_3:write_n
	wire  [31:0] mm_interconnect_0_hex_3_s1_writedata;                      // mm_interconnect_0:HEX_3_s1_writedata -> HEX_3:writedata
	wire         mm_interconnect_0_hex_4_s1_chipselect;                     // mm_interconnect_0:HEX_4_s1_chipselect -> HEX_4:chipselect
	wire  [31:0] mm_interconnect_0_hex_4_s1_readdata;                       // HEX_4:readdata -> mm_interconnect_0:HEX_4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_4_s1_address;                        // mm_interconnect_0:HEX_4_s1_address -> HEX_4:address
	wire         mm_interconnect_0_hex_4_s1_write;                          // mm_interconnect_0:HEX_4_s1_write -> HEX_4:write_n
	wire  [31:0] mm_interconnect_0_hex_4_s1_writedata;                      // mm_interconnect_0:HEX_4_s1_writedata -> HEX_4:writedata
	wire         mm_interconnect_0_hex_5_s1_chipselect;                     // mm_interconnect_0:HEX_5_s1_chipselect -> HEX_5:chipselect
	wire  [31:0] mm_interconnect_0_hex_5_s1_readdata;                       // HEX_5:readdata -> mm_interconnect_0:HEX_5_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_5_s1_address;                        // mm_interconnect_0:HEX_5_s1_address -> HEX_5:address
	wire         mm_interconnect_0_hex_5_s1_write;                          // mm_interconnect_0:HEX_5_s1_write -> HEX_5:write_n
	wire  [31:0] mm_interconnect_0_hex_5_s1_writedata;                      // mm_interconnect_0:HEX_5_s1_writedata -> HEX_5:writedata
	wire         mm_interconnect_0_led_s1_chipselect;                       // mm_interconnect_0:LED_s1_chipselect -> LED:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                         // LED:readdata -> mm_interconnect_0:LED_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                          // mm_interconnect_0:LED_s1_address -> LED:address
	wire         mm_interconnect_0_led_s1_write;                            // mm_interconnect_0:LED_s1_write -> LED:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                        // mm_interconnect_0:LED_s1_writedata -> LED:writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> CPU:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [CODE_MEMORY:reset, CPU:reset_n, HEX_0:reset_n, HEX_1:reset_n, HEX_2:reset_n, HEX_3:reset_n, HEX_4:reset_n, HEX_5:reset_n, LED:reset_n, TL_0:reset_n, TL_1:reset_n, TL_2:reset_n, TL_3:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sysid:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [CODE_MEMORY:reset_req, CPU:reset_req, rst_translator:reset_req_in]

	traffic_light_CODE_MEMORY code_memory (
		.clk        (clk_clk),                                     //   clk1.clk
		.address    (mm_interconnect_0_code_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_code_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_code_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_code_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_code_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_code_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_code_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze     (1'b0)                                         // (terminated)
	);

	traffic_light_CPU cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	traffic_light_HEX_0 hex_0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_0_s1_readdata),   //                    .readdata
		.out_port   (hex_0_external_connection_export)       // external_connection.export
	);

	traffic_light_HEX_0 hex_1 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_1_s1_readdata),   //                    .readdata
		.out_port   (hex_1_external_connection_export)       // external_connection.export
	);

	traffic_light_HEX_2 hex_2 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_2_s1_readdata),   //                    .readdata
		.out_port   (hex_2_external_connection_export)       // external_connection.export
	);

	traffic_light_HEX_2 hex_3 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_3_s1_readdata),   //                    .readdata
		.out_port   (hex_3_external_connection_export)       // external_connection.export
	);

	traffic_light_HEX_2 hex_4 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_4_s1_readdata),   //                    .readdata
		.out_port   (hex_4_external_connection_export)       // external_connection.export
	);

	traffic_light_HEX_2 hex_5 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hex_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_5_s1_readdata),   //                    .readdata
		.out_port   (hex_5_external_connection_export)       // external_connection.export
	);

	traffic_light_LED led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	traffic_light_TL_0 tl_0 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_tl_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tl_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tl_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tl_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tl_0_s1_readdata),   //                    .readdata
		.out_port   (tl_0_external_connection_export)       // external_connection.export
	);

	traffic_light_TL_0 tl_1 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_tl_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tl_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tl_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tl_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tl_1_s1_readdata),   //                    .readdata
		.out_port   (tl_1_external_connection_export)       // external_connection.export
	);

	traffic_light_TL_0 tl_2 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_tl_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tl_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tl_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tl_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tl_2_s1_readdata),   //                    .readdata
		.out_port   (tl_2_external_connection_export)       // external_connection.export
	);

	traffic_light_TL_0 tl_3 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_tl_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tl_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tl_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tl_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tl_3_s1_readdata),   //                    .readdata
		.out_port   (tl_3_external_connection_export)       // external_connection.export
	);

	traffic_light_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	traffic_light_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	traffic_light_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	traffic_light_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                           (clk_clk),                                                   //                       clk_0_clk.clk
		.CPU_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                            // CPU_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address                 (cpu_data_master_address),                                   //                 CPU_data_master.address
		.CPU_data_master_waitrequest             (cpu_data_master_waitrequest),                               //                                .waitrequest
		.CPU_data_master_byteenable              (cpu_data_master_byteenable),                                //                                .byteenable
		.CPU_data_master_read                    (cpu_data_master_read),                                      //                                .read
		.CPU_data_master_readdata                (cpu_data_master_readdata),                                  //                                .readdata
		.CPU_data_master_write                   (cpu_data_master_write),                                     //                                .write
		.CPU_data_master_writedata               (cpu_data_master_writedata),                                 //                                .writedata
		.CPU_data_master_debugaccess             (cpu_data_master_debugaccess),                               //                                .debugaccess
		.CPU_instruction_master_address          (cpu_instruction_master_address),                            //          CPU_instruction_master.address
		.CPU_instruction_master_waitrequest      (cpu_instruction_master_waitrequest),                        //                                .waitrequest
		.CPU_instruction_master_read             (cpu_instruction_master_read),                               //                                .read
		.CPU_instruction_master_readdata         (cpu_instruction_master_readdata),                           //                                .readdata
		.CODE_MEMORY_s1_address                  (mm_interconnect_0_code_memory_s1_address),                  //                  CODE_MEMORY_s1.address
		.CODE_MEMORY_s1_write                    (mm_interconnect_0_code_memory_s1_write),                    //                                .write
		.CODE_MEMORY_s1_readdata                 (mm_interconnect_0_code_memory_s1_readdata),                 //                                .readdata
		.CODE_MEMORY_s1_writedata                (mm_interconnect_0_code_memory_s1_writedata),                //                                .writedata
		.CODE_MEMORY_s1_byteenable               (mm_interconnect_0_code_memory_s1_byteenable),               //                                .byteenable
		.CODE_MEMORY_s1_chipselect               (mm_interconnect_0_code_memory_s1_chipselect),               //                                .chipselect
		.CODE_MEMORY_s1_clken                    (mm_interconnect_0_code_memory_s1_clken),                    //                                .clken
		.CPU_debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),             //             CPU_debug_mem_slave.address
		.CPU_debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                .write
		.CPU_debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                .read
		.CPU_debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                .readdata
		.CPU_debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                .writedata
		.CPU_debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                .byteenable
		.CPU_debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                .waitrequest
		.CPU_debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                .debugaccess
		.HEX_0_s1_address                        (mm_interconnect_0_hex_0_s1_address),                        //                        HEX_0_s1.address
		.HEX_0_s1_write                          (mm_interconnect_0_hex_0_s1_write),                          //                                .write
		.HEX_0_s1_readdata                       (mm_interconnect_0_hex_0_s1_readdata),                       //                                .readdata
		.HEX_0_s1_writedata                      (mm_interconnect_0_hex_0_s1_writedata),                      //                                .writedata
		.HEX_0_s1_chipselect                     (mm_interconnect_0_hex_0_s1_chipselect),                     //                                .chipselect
		.HEX_1_s1_address                        (mm_interconnect_0_hex_1_s1_address),                        //                        HEX_1_s1.address
		.HEX_1_s1_write                          (mm_interconnect_0_hex_1_s1_write),                          //                                .write
		.HEX_1_s1_readdata                       (mm_interconnect_0_hex_1_s1_readdata),                       //                                .readdata
		.HEX_1_s1_writedata                      (mm_interconnect_0_hex_1_s1_writedata),                      //                                .writedata
		.HEX_1_s1_chipselect                     (mm_interconnect_0_hex_1_s1_chipselect),                     //                                .chipselect
		.HEX_2_s1_address                        (mm_interconnect_0_hex_2_s1_address),                        //                        HEX_2_s1.address
		.HEX_2_s1_write                          (mm_interconnect_0_hex_2_s1_write),                          //                                .write
		.HEX_2_s1_readdata                       (mm_interconnect_0_hex_2_s1_readdata),                       //                                .readdata
		.HEX_2_s1_writedata                      (mm_interconnect_0_hex_2_s1_writedata),                      //                                .writedata
		.HEX_2_s1_chipselect                     (mm_interconnect_0_hex_2_s1_chipselect),                     //                                .chipselect
		.HEX_3_s1_address                        (mm_interconnect_0_hex_3_s1_address),                        //                        HEX_3_s1.address
		.HEX_3_s1_write                          (mm_interconnect_0_hex_3_s1_write),                          //                                .write
		.HEX_3_s1_readdata                       (mm_interconnect_0_hex_3_s1_readdata),                       //                                .readdata
		.HEX_3_s1_writedata                      (mm_interconnect_0_hex_3_s1_writedata),                      //                                .writedata
		.HEX_3_s1_chipselect                     (mm_interconnect_0_hex_3_s1_chipselect),                     //                                .chipselect
		.HEX_4_s1_address                        (mm_interconnect_0_hex_4_s1_address),                        //                        HEX_4_s1.address
		.HEX_4_s1_write                          (mm_interconnect_0_hex_4_s1_write),                          //                                .write
		.HEX_4_s1_readdata                       (mm_interconnect_0_hex_4_s1_readdata),                       //                                .readdata
		.HEX_4_s1_writedata                      (mm_interconnect_0_hex_4_s1_writedata),                      //                                .writedata
		.HEX_4_s1_chipselect                     (mm_interconnect_0_hex_4_s1_chipselect),                     //                                .chipselect
		.HEX_5_s1_address                        (mm_interconnect_0_hex_5_s1_address),                        //                        HEX_5_s1.address
		.HEX_5_s1_write                          (mm_interconnect_0_hex_5_s1_write),                          //                                .write
		.HEX_5_s1_readdata                       (mm_interconnect_0_hex_5_s1_readdata),                       //                                .readdata
		.HEX_5_s1_writedata                      (mm_interconnect_0_hex_5_s1_writedata),                      //                                .writedata
		.HEX_5_s1_chipselect                     (mm_interconnect_0_hex_5_s1_chipselect),                     //                                .chipselect
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                .chipselect
		.LED_s1_address                          (mm_interconnect_0_led_s1_address),                          //                          LED_s1.address
		.LED_s1_write                            (mm_interconnect_0_led_s1_write),                            //                                .write
		.LED_s1_readdata                         (mm_interconnect_0_led_s1_readdata),                         //                                .readdata
		.LED_s1_writedata                        (mm_interconnect_0_led_s1_writedata),                        //                                .writedata
		.LED_s1_chipselect                       (mm_interconnect_0_led_s1_chipselect),                       //                                .chipselect
		.sysid_control_slave_address             (mm_interconnect_0_sysid_control_slave_address),             //             sysid_control_slave.address
		.sysid_control_slave_readdata            (mm_interconnect_0_sysid_control_slave_readdata),            //                                .readdata
		.timer_0_s1_address                      (mm_interconnect_0_timer_0_s1_address),                      //                      timer_0_s1.address
		.timer_0_s1_write                        (mm_interconnect_0_timer_0_s1_write),                        //                                .write
		.timer_0_s1_readdata                     (mm_interconnect_0_timer_0_s1_readdata),                     //                                .readdata
		.timer_0_s1_writedata                    (mm_interconnect_0_timer_0_s1_writedata),                    //                                .writedata
		.timer_0_s1_chipselect                   (mm_interconnect_0_timer_0_s1_chipselect),                   //                                .chipselect
		.TL_0_s1_address                         (mm_interconnect_0_tl_0_s1_address),                         //                         TL_0_s1.address
		.TL_0_s1_write                           (mm_interconnect_0_tl_0_s1_write),                           //                                .write
		.TL_0_s1_readdata                        (mm_interconnect_0_tl_0_s1_readdata),                        //                                .readdata
		.TL_0_s1_writedata                       (mm_interconnect_0_tl_0_s1_writedata),                       //                                .writedata
		.TL_0_s1_chipselect                      (mm_interconnect_0_tl_0_s1_chipselect),                      //                                .chipselect
		.TL_1_s1_address                         (mm_interconnect_0_tl_1_s1_address),                         //                         TL_1_s1.address
		.TL_1_s1_write                           (mm_interconnect_0_tl_1_s1_write),                           //                                .write
		.TL_1_s1_readdata                        (mm_interconnect_0_tl_1_s1_readdata),                        //                                .readdata
		.TL_1_s1_writedata                       (mm_interconnect_0_tl_1_s1_writedata),                       //                                .writedata
		.TL_1_s1_chipselect                      (mm_interconnect_0_tl_1_s1_chipselect),                      //                                .chipselect
		.TL_2_s1_address                         (mm_interconnect_0_tl_2_s1_address),                         //                         TL_2_s1.address
		.TL_2_s1_write                           (mm_interconnect_0_tl_2_s1_write),                           //                                .write
		.TL_2_s1_readdata                        (mm_interconnect_0_tl_2_s1_readdata),                        //                                .readdata
		.TL_2_s1_writedata                       (mm_interconnect_0_tl_2_s1_writedata),                       //                                .writedata
		.TL_2_s1_chipselect                      (mm_interconnect_0_tl_2_s1_chipselect),                      //                                .chipselect
		.TL_3_s1_address                         (mm_interconnect_0_tl_3_s1_address),                         //                         TL_3_s1.address
		.TL_3_s1_write                           (mm_interconnect_0_tl_3_s1_write),                           //                                .write
		.TL_3_s1_readdata                        (mm_interconnect_0_tl_3_s1_readdata),                        //                                .readdata
		.TL_3_s1_writedata                       (mm_interconnect_0_tl_3_s1_writedata),                       //                                .writedata
		.TL_3_s1_chipselect                      (mm_interconnect_0_tl_3_s1_chipselect)                       //                                .chipselect
	);

	traffic_light_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
